package NbiFullAdder;


(*synthesize*)
module mkNbFA()

endpackage: NbiFullAdder
